library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

package matrix_pkg is
    -- ????
    type STD_LOGIC_VECTOR_ARRAY is array (0 to 127) of STD_LOGIC_VECTOR(7 downto 0);
end package matrix_pkg;
