library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package config_pkg is
    constant WIDTH : integer := 256;  -- ????
end package config_pkg;

